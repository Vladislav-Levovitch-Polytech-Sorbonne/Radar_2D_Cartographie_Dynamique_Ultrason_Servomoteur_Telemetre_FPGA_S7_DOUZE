
module Neopixel (
	clk_clk,
	reset_reset_n,
	neopixel_alone_output_commande_neopixel);	

	input		clk_clk;
	input		reset_reset_n;
	output		neopixel_alone_output_commande_neopixel;
endmodule
