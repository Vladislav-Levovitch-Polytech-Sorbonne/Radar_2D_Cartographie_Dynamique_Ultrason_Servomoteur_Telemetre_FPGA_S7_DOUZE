
module Neopixel_Alone_bis (
	clk_clk,
	neopixel_alone_output_commande_neopixel,
	reset_reset_n);	

	input		clk_clk;
	output		neopixel_alone_output_commande_neopixel;
	input		reset_reset_n;
endmodule
