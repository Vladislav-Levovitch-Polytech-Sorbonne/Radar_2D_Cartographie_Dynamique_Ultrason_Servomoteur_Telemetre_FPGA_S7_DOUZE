// Neopixel_Neopixel_0.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module Neopixel_Neopixel_0 (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	Neopixel_Neopixel_0_Neopixel_0 neopixel_0 (
	);

endmodule
